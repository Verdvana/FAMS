// qsys_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module qsys_system (
		input  wire [23:0] adc_p_export,      //      adc_p.export
		input  wire [23:0] adc_t_export,      //      adc_t.export
		input  wire        clk_clk,           //        clk.clk
		input  wire [15:0] dig_p1_export,     //     dig_p1.export
		input  wire [15:0] dig_p2_export,     //     dig_p2.export
		input  wire [15:0] dig_p3_export,     //     dig_p3.export
		input  wire [15:0] dig_p4_export,     //     dig_p4.export
		input  wire [15:0] dig_p5_export,     //     dig_p5.export
		input  wire [15:0] dig_p6_export,     //     dig_p6.export
		input  wire [15:0] dig_p7_export,     //     dig_p7.export
		input  wire [15:0] dig_p8_export,     //     dig_p8.export
		input  wire [15:0] dig_p9_export,     //     dig_p9.export
		input  wire [15:0] dig_t1_export,     //     dig_t1.export
		input  wire [15:0] dig_t2_export,     //     dig_t2.export
		input  wire [15:0] dig_t3_export,     //     dig_t3.export
		input  wire        end_o_export,      //      end_o.export
		output wire [7:0]  heart_rate_export, // heart_rate.export
		output wire [7:0]  heignt_dec_export, // heignt_dec.export
		output wire [7:0]  heignt_int_export, // heignt_int.export
		input  wire [23:0] max30102_0_export, // max30102_0.export
		input  wire [23:0] max30102_1_export, // max30102_1.export
		input  wire        reset_reset_n      //      reset.reset_n
	);

	wire  [31:0] nios2_gen2_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire         nios2_gen2_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire         nios2_gen2_data_master_debugaccess;                        // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	wire  [16:0] nios2_gen2_data_master_address;                            // nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	wire   [3:0] nios2_gen2_data_master_byteenable;                         // nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	wire         nios2_gen2_data_master_read;                               // nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	wire         nios2_gen2_data_master_readdatavalid;                      // mm_interconnect_0:nios2_gen2_data_master_readdatavalid -> nios2_gen2:d_readdatavalid
	wire         nios2_gen2_data_master_write;                              // nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	wire  [31:0] nios2_gen2_data_master_writedata;                          // nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	wire  [31:0] nios2_gen2_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire         nios2_gen2_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire  [16:0] nios2_gen2_instruction_master_address;                     // nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	wire         nios2_gen2_instruction_master_read;                        // nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	wire         nios2_gen2_instruction_master_readdatavalid;               // mm_interconnect_0:nios2_gen2_instruction_master_readdatavalid -> nios2_gen2:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;       // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;        // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata;     // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest;  // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                       // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                         // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [12:0] mm_interconnect_0_ram_s1_address;                          // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                       // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                            // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                        // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                            // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire  [31:0] mm_interconnect_0_max30102_0_s1_readdata;                  // max30102_0:readdata -> mm_interconnect_0:max30102_0_s1_readdata
	wire   [1:0] mm_interconnect_0_max30102_0_s1_address;                   // mm_interconnect_0:max30102_0_s1_address -> max30102_0:address
	wire  [31:0] mm_interconnect_0_max30102_1_s1_readdata;                  // max30102_1:readdata -> mm_interconnect_0:max30102_1_s1_readdata
	wire   [1:0] mm_interconnect_0_max30102_1_s1_address;                   // mm_interconnect_0:max30102_1_s1_address -> max30102_1:address
	wire  [31:0] mm_interconnect_0_end_o_s1_readdata;                       // end_o:readdata -> mm_interconnect_0:end_o_s1_readdata
	wire   [1:0] mm_interconnect_0_end_o_s1_address;                        // mm_interconnect_0:end_o_s1_address -> end_o:address
	wire         mm_interconnect_0_heignt_int_s1_chipselect;                // mm_interconnect_0:heignt_int_s1_chipselect -> heignt_int:chipselect
	wire  [31:0] mm_interconnect_0_heignt_int_s1_readdata;                  // heignt_int:readdata -> mm_interconnect_0:heignt_int_s1_readdata
	wire   [1:0] mm_interconnect_0_heignt_int_s1_address;                   // mm_interconnect_0:heignt_int_s1_address -> heignt_int:address
	wire         mm_interconnect_0_heignt_int_s1_write;                     // mm_interconnect_0:heignt_int_s1_write -> heignt_int:write_n
	wire  [31:0] mm_interconnect_0_heignt_int_s1_writedata;                 // mm_interconnect_0:heignt_int_s1_writedata -> heignt_int:writedata
	wire         mm_interconnect_0_heignt_dec_s1_chipselect;                // mm_interconnect_0:heignt_dec_s1_chipselect -> heignt_dec:chipselect
	wire  [31:0] mm_interconnect_0_heignt_dec_s1_readdata;                  // heignt_dec:readdata -> mm_interconnect_0:heignt_dec_s1_readdata
	wire   [1:0] mm_interconnect_0_heignt_dec_s1_address;                   // mm_interconnect_0:heignt_dec_s1_address -> heignt_dec:address
	wire         mm_interconnect_0_heignt_dec_s1_write;                     // mm_interconnect_0:heignt_dec_s1_write -> heignt_dec:write_n
	wire  [31:0] mm_interconnect_0_heignt_dec_s1_writedata;                 // mm_interconnect_0:heignt_dec_s1_writedata -> heignt_dec:writedata
	wire         mm_interconnect_0_heart_rate_s1_chipselect;                // mm_interconnect_0:heart_rate_s1_chipselect -> heart_rate:chipselect
	wire  [31:0] mm_interconnect_0_heart_rate_s1_readdata;                  // heart_rate:readdata -> mm_interconnect_0:heart_rate_s1_readdata
	wire   [1:0] mm_interconnect_0_heart_rate_s1_address;                   // mm_interconnect_0:heart_rate_s1_address -> heart_rate:address
	wire         mm_interconnect_0_heart_rate_s1_write;                     // mm_interconnect_0:heart_rate_s1_write -> heart_rate:write_n
	wire  [31:0] mm_interconnect_0_heart_rate_s1_writedata;                 // mm_interconnect_0:heart_rate_s1_writedata -> heart_rate:writedata
	wire  [31:0] mm_interconnect_0_dig_t1_s1_readdata;                      // dig_t1:readdata -> mm_interconnect_0:dig_t1_s1_readdata
	wire   [1:0] mm_interconnect_0_dig_t1_s1_address;                       // mm_interconnect_0:dig_t1_s1_address -> dig_t1:address
	wire  [31:0] mm_interconnect_0_dig_t2_s1_readdata;                      // dig_t2:readdata -> mm_interconnect_0:dig_t2_s1_readdata
	wire   [1:0] mm_interconnect_0_dig_t2_s1_address;                       // mm_interconnect_0:dig_t2_s1_address -> dig_t2:address
	wire  [31:0] mm_interconnect_0_dig_t3_s1_readdata;                      // dig_t3:readdata -> mm_interconnect_0:dig_t3_s1_readdata
	wire   [1:0] mm_interconnect_0_dig_t3_s1_address;                       // mm_interconnect_0:dig_t3_s1_address -> dig_t3:address
	wire  [31:0] mm_interconnect_0_dig_p1_s1_readdata;                      // dig_p1:readdata -> mm_interconnect_0:dig_p1_s1_readdata
	wire   [1:0] mm_interconnect_0_dig_p1_s1_address;                       // mm_interconnect_0:dig_p1_s1_address -> dig_p1:address
	wire  [31:0] mm_interconnect_0_dig_p2_s1_readdata;                      // dig_p2:readdata -> mm_interconnect_0:dig_p2_s1_readdata
	wire   [1:0] mm_interconnect_0_dig_p2_s1_address;                       // mm_interconnect_0:dig_p2_s1_address -> dig_p2:address
	wire  [31:0] mm_interconnect_0_dig_p3_s1_readdata;                      // dig_p3:readdata -> mm_interconnect_0:dig_p3_s1_readdata
	wire   [1:0] mm_interconnect_0_dig_p3_s1_address;                       // mm_interconnect_0:dig_p3_s1_address -> dig_p3:address
	wire  [31:0] mm_interconnect_0_dig_p4_s1_readdata;                      // dig_p4:readdata -> mm_interconnect_0:dig_p4_s1_readdata
	wire   [1:0] mm_interconnect_0_dig_p4_s1_address;                       // mm_interconnect_0:dig_p4_s1_address -> dig_p4:address
	wire  [31:0] mm_interconnect_0_dig_p6_s1_readdata;                      // dig_p6:readdata -> mm_interconnect_0:dig_p6_s1_readdata
	wire   [1:0] mm_interconnect_0_dig_p6_s1_address;                       // mm_interconnect_0:dig_p6_s1_address -> dig_p6:address
	wire  [31:0] mm_interconnect_0_dig_p5_s1_readdata;                      // dig_p5:readdata -> mm_interconnect_0:dig_p5_s1_readdata
	wire   [1:0] mm_interconnect_0_dig_p5_s1_address;                       // mm_interconnect_0:dig_p5_s1_address -> dig_p5:address
	wire  [31:0] mm_interconnect_0_dig_p7_s1_readdata;                      // dig_p7:readdata -> mm_interconnect_0:dig_p7_s1_readdata
	wire   [1:0] mm_interconnect_0_dig_p7_s1_address;                       // mm_interconnect_0:dig_p7_s1_address -> dig_p7:address
	wire  [31:0] mm_interconnect_0_dig_p8_s1_readdata;                      // dig_p8:readdata -> mm_interconnect_0:dig_p8_s1_readdata
	wire   [1:0] mm_interconnect_0_dig_p8_s1_address;                       // mm_interconnect_0:dig_p8_s1_address -> dig_p8:address
	wire  [31:0] mm_interconnect_0_dig_p9_s1_readdata;                      // dig_p9:readdata -> mm_interconnect_0:dig_p9_s1_readdata
	wire   [1:0] mm_interconnect_0_dig_p9_s1_address;                       // mm_interconnect_0:dig_p9_s1_address -> dig_p9:address
	wire  [31:0] mm_interconnect_0_adc_t_s1_readdata;                       // adc_t:readdata -> mm_interconnect_0:adc_t_s1_readdata
	wire   [1:0] mm_interconnect_0_adc_t_s1_address;                        // mm_interconnect_0:adc_t_s1_address -> adc_t:address
	wire  [31:0] mm_interconnect_0_adc_p_s1_readdata;                       // adc_p:readdata -> mm_interconnect_0:adc_p_s1_readdata
	wire   [1:0] mm_interconnect_0_adc_p_s1_address;                        // mm_interconnect_0:adc_p_s1_address -> adc_p:address
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [RAM:reset, adc_p:reset_n, adc_t:reset_n, dig_p1:reset_n, dig_p2:reset_n, dig_p3:reset_n, dig_p4:reset_n, dig_p5:reset_n, dig_p6:reset_n, dig_p7:reset_n, dig_p8:reset_n, dig_p9:reset_n, dig_t1:reset_n, dig_t2:reset_n, dig_t3:reset_n, end_o:reset_n, heart_rate:reset_n, heignt_dec:reset_n, heignt_int:reset_n, irq_mapper:reset, jtag_uart:rst_n, max30102_0:reset_n, max30102_1:reset_n, mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n, rst_translator:in_reset, sysid_qsys:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [RAM:reset_req, nios2_gen2:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_debug_reset_request_reset;                      // nios2_gen2:debug_reset_request -> rst_controller:reset_in1

	qsys_system_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	qsys_system_adc_p adc_p (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_adc_p_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_adc_p_s1_readdata), //                    .readdata
		.in_port  (adc_p_export)                         // external_connection.export
	);

	qsys_system_adc_p adc_t (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_adc_t_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_adc_t_s1_readdata), //                    .readdata
		.in_port  (adc_t_export)                         // external_connection.export
	);

	qsys_system_dig_p1 dig_p1 (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_dig_p1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dig_p1_s1_readdata), //                    .readdata
		.in_port  (dig_p1_export)                         // external_connection.export
	);

	qsys_system_dig_p1 dig_p2 (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_dig_p2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dig_p2_s1_readdata), //                    .readdata
		.in_port  (dig_p2_export)                         // external_connection.export
	);

	qsys_system_dig_p1 dig_p3 (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_dig_p3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dig_p3_s1_readdata), //                    .readdata
		.in_port  (dig_p3_export)                         // external_connection.export
	);

	qsys_system_dig_p1 dig_p4 (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_dig_p4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dig_p4_s1_readdata), //                    .readdata
		.in_port  (dig_p4_export)                         // external_connection.export
	);

	qsys_system_dig_p1 dig_p5 (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_dig_p5_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dig_p5_s1_readdata), //                    .readdata
		.in_port  (dig_p5_export)                         // external_connection.export
	);

	qsys_system_dig_p1 dig_p6 (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_dig_p6_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dig_p6_s1_readdata), //                    .readdata
		.in_port  (dig_p6_export)                         // external_connection.export
	);

	qsys_system_dig_p1 dig_p7 (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_dig_p7_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dig_p7_s1_readdata), //                    .readdata
		.in_port  (dig_p7_export)                         // external_connection.export
	);

	qsys_system_dig_p1 dig_p8 (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_dig_p8_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dig_p8_s1_readdata), //                    .readdata
		.in_port  (dig_p8_export)                         // external_connection.export
	);

	qsys_system_dig_p1 dig_p9 (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_dig_p9_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dig_p9_s1_readdata), //                    .readdata
		.in_port  (dig_p9_export)                         // external_connection.export
	);

	qsys_system_dig_p1 dig_t1 (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_dig_t1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dig_t1_s1_readdata), //                    .readdata
		.in_port  (dig_t1_export)                         // external_connection.export
	);

	qsys_system_dig_p1 dig_t2 (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_dig_t2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dig_t2_s1_readdata), //                    .readdata
		.in_port  (dig_t2_export)                         // external_connection.export
	);

	qsys_system_dig_p1 dig_t3 (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_dig_t3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dig_t3_s1_readdata), //                    .readdata
		.in_port  (dig_t3_export)                         // external_connection.export
	);

	qsys_system_end_o end_o (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_end_o_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_end_o_s1_readdata), //                    .readdata
		.in_port  (end_o_export)                         // external_connection.export
	);

	qsys_system_heart_rate heart_rate (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_heart_rate_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_heart_rate_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_heart_rate_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_heart_rate_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_heart_rate_s1_readdata),   //                    .readdata
		.out_port   (heart_rate_export)                           // external_connection.export
	);

	qsys_system_heart_rate heignt_dec (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_heignt_dec_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_heignt_dec_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_heignt_dec_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_heignt_dec_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_heignt_dec_s1_readdata),   //                    .readdata
		.out_port   (heignt_dec_export)                           // external_connection.export
	);

	qsys_system_heart_rate heignt_int (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_heignt_int_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_heignt_int_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_heignt_int_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_heignt_int_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_heignt_int_s1_readdata),   //                    .readdata
		.out_port   (heignt_int_export)                           // external_connection.export
	);

	qsys_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	qsys_system_adc_p max30102_0 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_max30102_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_max30102_0_s1_readdata), //                    .readdata
		.in_port  (max30102_0_export)                         // external_connection.export
	);

	qsys_system_adc_p max30102_1 (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_max30102_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_max30102_1_s1_readdata), //                    .readdata
		.in_port  (max30102_1_export)                         // external_connection.export
	);

	qsys_system_nios2_gen2 nios2_gen2 (
		.clk                                 (clk_clk),                                                  //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                          //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                       //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	qsys_system_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	qsys_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                  (clk_clk),                                                   //                                clk_clk.clk
		.nios2_gen2_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // nios2_gen2_reset_reset_bridge_in_reset.reset
		.nios2_gen2_data_master_address               (nios2_gen2_data_master_address),                            //                 nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest           (nios2_gen2_data_master_waitrequest),                        //                                       .waitrequest
		.nios2_gen2_data_master_byteenable            (nios2_gen2_data_master_byteenable),                         //                                       .byteenable
		.nios2_gen2_data_master_read                  (nios2_gen2_data_master_read),                               //                                       .read
		.nios2_gen2_data_master_readdata              (nios2_gen2_data_master_readdata),                           //                                       .readdata
		.nios2_gen2_data_master_readdatavalid         (nios2_gen2_data_master_readdatavalid),                      //                                       .readdatavalid
		.nios2_gen2_data_master_write                 (nios2_gen2_data_master_write),                              //                                       .write
		.nios2_gen2_data_master_writedata             (nios2_gen2_data_master_writedata),                          //                                       .writedata
		.nios2_gen2_data_master_debugaccess           (nios2_gen2_data_master_debugaccess),                        //                                       .debugaccess
		.nios2_gen2_instruction_master_address        (nios2_gen2_instruction_master_address),                     //          nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest    (nios2_gen2_instruction_master_waitrequest),                 //                                       .waitrequest
		.nios2_gen2_instruction_master_read           (nios2_gen2_instruction_master_read),                        //                                       .read
		.nios2_gen2_instruction_master_readdata       (nios2_gen2_instruction_master_readdata),                    //                                       .readdata
		.nios2_gen2_instruction_master_readdatavalid  (nios2_gen2_instruction_master_readdatavalid),               //                                       .readdatavalid
		.adc_p_s1_address                             (mm_interconnect_0_adc_p_s1_address),                        //                               adc_p_s1.address
		.adc_p_s1_readdata                            (mm_interconnect_0_adc_p_s1_readdata),                       //                                       .readdata
		.adc_t_s1_address                             (mm_interconnect_0_adc_t_s1_address),                        //                               adc_t_s1.address
		.adc_t_s1_readdata                            (mm_interconnect_0_adc_t_s1_readdata),                       //                                       .readdata
		.dig_p1_s1_address                            (mm_interconnect_0_dig_p1_s1_address),                       //                              dig_p1_s1.address
		.dig_p1_s1_readdata                           (mm_interconnect_0_dig_p1_s1_readdata),                      //                                       .readdata
		.dig_p2_s1_address                            (mm_interconnect_0_dig_p2_s1_address),                       //                              dig_p2_s1.address
		.dig_p2_s1_readdata                           (mm_interconnect_0_dig_p2_s1_readdata),                      //                                       .readdata
		.dig_p3_s1_address                            (mm_interconnect_0_dig_p3_s1_address),                       //                              dig_p3_s1.address
		.dig_p3_s1_readdata                           (mm_interconnect_0_dig_p3_s1_readdata),                      //                                       .readdata
		.dig_p4_s1_address                            (mm_interconnect_0_dig_p4_s1_address),                       //                              dig_p4_s1.address
		.dig_p4_s1_readdata                           (mm_interconnect_0_dig_p4_s1_readdata),                      //                                       .readdata
		.dig_p5_s1_address                            (mm_interconnect_0_dig_p5_s1_address),                       //                              dig_p5_s1.address
		.dig_p5_s1_readdata                           (mm_interconnect_0_dig_p5_s1_readdata),                      //                                       .readdata
		.dig_p6_s1_address                            (mm_interconnect_0_dig_p6_s1_address),                       //                              dig_p6_s1.address
		.dig_p6_s1_readdata                           (mm_interconnect_0_dig_p6_s1_readdata),                      //                                       .readdata
		.dig_p7_s1_address                            (mm_interconnect_0_dig_p7_s1_address),                       //                              dig_p7_s1.address
		.dig_p7_s1_readdata                           (mm_interconnect_0_dig_p7_s1_readdata),                      //                                       .readdata
		.dig_p8_s1_address                            (mm_interconnect_0_dig_p8_s1_address),                       //                              dig_p8_s1.address
		.dig_p8_s1_readdata                           (mm_interconnect_0_dig_p8_s1_readdata),                      //                                       .readdata
		.dig_p9_s1_address                            (mm_interconnect_0_dig_p9_s1_address),                       //                              dig_p9_s1.address
		.dig_p9_s1_readdata                           (mm_interconnect_0_dig_p9_s1_readdata),                      //                                       .readdata
		.dig_t1_s1_address                            (mm_interconnect_0_dig_t1_s1_address),                       //                              dig_t1_s1.address
		.dig_t1_s1_readdata                           (mm_interconnect_0_dig_t1_s1_readdata),                      //                                       .readdata
		.dig_t2_s1_address                            (mm_interconnect_0_dig_t2_s1_address),                       //                              dig_t2_s1.address
		.dig_t2_s1_readdata                           (mm_interconnect_0_dig_t2_s1_readdata),                      //                                       .readdata
		.dig_t3_s1_address                            (mm_interconnect_0_dig_t3_s1_address),                       //                              dig_t3_s1.address
		.dig_t3_s1_readdata                           (mm_interconnect_0_dig_t3_s1_readdata),                      //                                       .readdata
		.end_o_s1_address                             (mm_interconnect_0_end_o_s1_address),                        //                               end_o_s1.address
		.end_o_s1_readdata                            (mm_interconnect_0_end_o_s1_readdata),                       //                                       .readdata
		.heart_rate_s1_address                        (mm_interconnect_0_heart_rate_s1_address),                   //                          heart_rate_s1.address
		.heart_rate_s1_write                          (mm_interconnect_0_heart_rate_s1_write),                     //                                       .write
		.heart_rate_s1_readdata                       (mm_interconnect_0_heart_rate_s1_readdata),                  //                                       .readdata
		.heart_rate_s1_writedata                      (mm_interconnect_0_heart_rate_s1_writedata),                 //                                       .writedata
		.heart_rate_s1_chipselect                     (mm_interconnect_0_heart_rate_s1_chipselect),                //                                       .chipselect
		.heignt_dec_s1_address                        (mm_interconnect_0_heignt_dec_s1_address),                   //                          heignt_dec_s1.address
		.heignt_dec_s1_write                          (mm_interconnect_0_heignt_dec_s1_write),                     //                                       .write
		.heignt_dec_s1_readdata                       (mm_interconnect_0_heignt_dec_s1_readdata),                  //                                       .readdata
		.heignt_dec_s1_writedata                      (mm_interconnect_0_heignt_dec_s1_writedata),                 //                                       .writedata
		.heignt_dec_s1_chipselect                     (mm_interconnect_0_heignt_dec_s1_chipselect),                //                                       .chipselect
		.heignt_int_s1_address                        (mm_interconnect_0_heignt_int_s1_address),                   //                          heignt_int_s1.address
		.heignt_int_s1_write                          (mm_interconnect_0_heignt_int_s1_write),                     //                                       .write
		.heignt_int_s1_readdata                       (mm_interconnect_0_heignt_int_s1_readdata),                  //                                       .readdata
		.heignt_int_s1_writedata                      (mm_interconnect_0_heignt_int_s1_writedata),                 //                                       .writedata
		.heignt_int_s1_chipselect                     (mm_interconnect_0_heignt_int_s1_chipselect),                //                                       .chipselect
		.jtag_uart_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                       .write
		.jtag_uart_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                       .read
		.jtag_uart_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                       .chipselect
		.max30102_0_s1_address                        (mm_interconnect_0_max30102_0_s1_address),                   //                          max30102_0_s1.address
		.max30102_0_s1_readdata                       (mm_interconnect_0_max30102_0_s1_readdata),                  //                                       .readdata
		.max30102_1_s1_address                        (mm_interconnect_0_max30102_1_s1_address),                   //                          max30102_1_s1.address
		.max30102_1_s1_readdata                       (mm_interconnect_0_max30102_1_s1_readdata),                  //                                       .readdata
		.nios2_gen2_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),      //             nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),        //                                       .write
		.nios2_gen2_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),         //                                       .read
		.nios2_gen2_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),     //                                       .readdata
		.nios2_gen2_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),    //                                       .writedata
		.nios2_gen2_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),   //                                       .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest),  //                                       .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess),  //                                       .debugaccess
		.RAM_s1_address                               (mm_interconnect_0_ram_s1_address),                          //                                 RAM_s1.address
		.RAM_s1_write                                 (mm_interconnect_0_ram_s1_write),                            //                                       .write
		.RAM_s1_readdata                              (mm_interconnect_0_ram_s1_readdata),                         //                                       .readdata
		.RAM_s1_writedata                             (mm_interconnect_0_ram_s1_writedata),                        //                                       .writedata
		.RAM_s1_byteenable                            (mm_interconnect_0_ram_s1_byteenable),                       //                                       .byteenable
		.RAM_s1_chipselect                            (mm_interconnect_0_ram_s1_chipselect),                       //                                       .chipselect
		.RAM_s1_clken                                 (mm_interconnect_0_ram_s1_clken),                            //                                       .clken
		.sysid_qsys_control_slave_address             (mm_interconnect_0_sysid_qsys_control_slave_address),        //               sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata            (mm_interconnect_0_sysid_qsys_control_slave_readdata)        //                                       .readdata
	);

	qsys_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_irq_irq)              //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),       // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),   //          .reset_req
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

endmodule
