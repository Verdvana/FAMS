module ROM_rh(
		input	[11:0]	address,
		input		clock,
		output  reg q 
		
);

always@(posedge clock)
begin
	case(address)
	8'd0 :   q=0;
	8'd1 :   q=0;
	8'd2 :   q=0;
	8'd3 :   q=0;
	8'd4 :   q=0;
	8'd5 :   q=0;
	8'd6 :   q=0;
	8'd7 :   q=0;
	8'd8 :   q=0;
	8'd9 :   q=0;
	8'd10 :  q=0;
	8'd11 :  q=0;
	8'd12 :  q=0;
	8'd13 :  q=0;
	8'd14 :  q=0;
	8'd15 :  q=0;
	8'd16 :  q=0;
	8'd17 :  q=0;
	8'd18 :  q=0;
	8'd19 :  q=0;
	8'd20 :  q=0;
	8'd21 :  q=0;
	8'd22 :  q=0;
	8'd23 :  q=0;
	8'd24 :  q=0;
	8'd25 :  q=0;
	8'd26 :  q=0;
	8'd27 :  q=0;
	8'd28 :  q=0;
	8'd29 :  q=0;
	8'd30 :  q=0;
	8'd31 :  q=0;
	8'd32 :  q=0;
	8'd33 :  q=0;
	8'd34 :  q=0;
	8'd35 :  q=0;
	8'd36 :  q=0;
	8'd37 :  q=0;
	8'd38 :  q=0;
	8'd39 :  q=0;
	8'd40 :  q=0;
	8'd41 :  q=0;
	8'd42 :  q=0;
	8'd43 :  q=0;
	8'd44 :  q=0;
	8'd45 :  q=0;
	8'd46 :  q=0;
	8'd47 :  q=0;
	8'd48 :  q=0;
	8'd49 :  q=1;
	8'd50 :  q=1;
	8'd51 :  q=1;
	8'd52 :  q=1;
	8'd53 :  q=1;
	8'd54 :  q=0;
	8'd55 :  q=0;
	8'd56 :  q=0;
	8'd57 :  q=1;
	8'd58 :  q=0;
	8'd59 :  q=0;
	8'd60 :  q=0;
	8'd61 :  q=0;
	8'd62 :  q=1;
	8'd63 :  q=0;
	8'd64 :  q=0;
	8'd65 :  q=1;
	8'd66 :  q=0;
	8'd67 :  q=0;
	8'd68 :  q=0;
	8'd69 :  q=1;
	8'd70 :  q=1;
	8'd71 :  q=0;
	8'd72 :  q=0;
	8'd73 :  q=1;
	8'd74 :  q=0;
	8'd75 :  q=0;
	8'd76 :  q=0;
	8'd77 :  q=0;
	8'd78 :  q=1;
	8'd79 :  q=0;
	8'd80 :  q=0;
	8'd81 :  q=1;
	8'd82 :  q=0;
	8'd83 :  q=0;
	8'd84 :  q=0;
	8'd85 :  q=0;
	8'd86 :  q=1;
	8'd87 :  q=0;
	8'd88 :  q=0;
	8'd89 :  q=1;
	8'd90 :  q=0;
	8'd91 :  q=0;
	8'd92 :  q=0;
	8'd93 :  q=0;
	8'd94 :  q=1;
	8'd95 :  q=0;
	8'd96 :  q=0;
	8'd97 :  q=1;
	8'd98 :  q=0;
	8'd99 :  q=0;
	8'd100 : q=0;
	8'd101 : q=0;
	8'd102 : q=1;
	8'd103 : q=0;
	8'd104 : q=0;
	8'd105 : q=1;
	8'd106 : q=0;
	8'd107 : q=0;
	8'd108 : q=0;
	8'd109 : q=0;
	8'd110 : q=1;
	8'd111 : q=0;
	8'd112 : q=0;
	8'd113 : q=1;
	8'd114 : q=0;
	8'd115 : q=0;
	8'd116 : q=0;
	8'd117 : q=1;
	8'd118 : q=1;
	8'd119 : q=0;
	8'd120 : q=0;
	8'd121 : q=1;
	8'd122 : q=1;
	8'd123 : q=1;
	8'd124 : q=1;
	8'd125 : q=1;
	8'd126 : q=1;
	8'd127 : q=0;
	8'd128 : q=0;
	8'd129 : q=1;
	8'd130 : q=1;
	8'd131 : q=1;
	8'd132 : q=1;
	8'd133 : q=1;
	8'd134 : q=0;
	8'd135 : q=0;
	8'd136 : q=0;
	8'd137 : q=1;
	8'd138 : q=1;
	8'd139 : q=1;
	8'd140 : q=1;
	8'd141 : q=1;
	8'd142 : q=1;
	8'd143 : q=0;
	8'd144 : q=0;
	8'd145 : q=1;
	8'd146 : q=0;
	8'd147 : q=0;
	8'd148 : q=1;
	8'd149 : q=0;
	8'd150 : q=0;
	8'd151 : q=0;
	8'd152 : q=0;
	8'd153 : q=1;
	8'd154 : q=0;
	8'd155 : q=0;
	8'd156 : q=0;
	8'd157 : q=0;
	8'd158 : q=1;
	8'd159 : q=0;
	8'd160 : q=0;
	8'd161 : q=1;
	8'd162 : q=0;
	8'd163 : q=0;
	8'd164 : q=1;
	8'd165 : q=1;
	8'd166 : q=0;
	8'd167 : q=0;
	8'd168 : q=0;
	8'd169 : q=1;
	8'd170 : q=0;
	8'd171 : q=0;
	8'd172 : q=0;
	8'd173 : q=0;
	8'd174 : q=1;
	8'd175 : q=0;
	8'd176 : q=0;
	8'd177 : q=1;
	8'd178 : q=0;
	8'd179 : q=0;
	8'd180 : q=0;
	8'd181 : q=1;
	8'd182 : q=0;
	8'd183 : q=0;
	8'd184 : q=0;
	8'd185 : q=1;
	8'd186 : q=0;
	8'd187 : q=0;
	8'd188 : q=0;
	8'd189 : q=0;
	8'd190 : q=1;
	8'd191 : q=0;
	8'd192 : q=0;
	8'd193 : q=1;
	8'd194 : q=0;
	8'd195 : q=0;
	8'd196 : q=0;
	8'd197 : q=1;
	8'd198 : q=1;
	8'd199 : q=0;
	8'd200 : q=0;
	8'd201 : q=1;
	8'd202 : q=0;
	8'd203 : q=0;
	8'd204 : q=0;
	8'd205 : q=0;
	8'd206 : q=1;
	8'd207 : q=0;
	8'd208 : q=0;
	8'd209 : q=1;
	8'd210 : q=0;
	8'd211 : q=0;
	8'd212 : q=0;
	8'd213 : q=0;
	8'd214 : q=1;
	8'd215 : q=0;
	8'd216 : q=0;
	8'd217 : q=1;
	8'd218 : q=0;
	8'd219 : q=0;
	8'd220 : q=0;
	8'd221 : q=0;
	8'd222 : q=1;
	8'd223 : q=0;
	8'd224 : q=0;
	8'd225 : q=0;
	8'd226 : q=0;
	8'd227 : q=0;
	8'd228 : q=0;
	8'd229 : q=0;
	8'd230 : q=0;
	8'd231 : q=0;
	8'd232 : q=0;
	8'd233 : q=0;
	8'd234 : q=0;
	8'd235 : q=0;
	8'd236 : q=0;
	8'd237 : q=0;
	8'd238 : q=0;
	8'd239 : q=0;
	8'd240 : q=0;
	8'd241 : q=0;
	8'd242 : q=0;
	8'd243 : q=0;
	8'd244 : q=0;
	8'd245 : q=0;
	8'd246 : q=0;
	8'd247 : q=0;
	8'd248 : q=0;
	8'd249 : q=0;
	8'd250 : q=0;
	8'd251 : q=0;
	8'd252 : q=0;
	8'd253 : q=0;
	8'd254 : q=0;
	8'd255 : q=0;		
		
	endcase
end




endmodule
